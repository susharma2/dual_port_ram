package pkg_b;

`include "define_file.sv"
`include "port_b_trans.sv"
`include "port_b_driver.sv"
`include "port_b_monitor.sv"

endpackage
