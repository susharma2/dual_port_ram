package pkg;

import pkg_a::*;
import pkg_b::*;

`include "define_file.sv"
`include "generator.sv"
`include "environment.sv"
`include "test.sv"

endpackage
