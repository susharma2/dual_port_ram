package pkg_a;

`include "define_file.sv"
`include "port_a_trans.sv"
`include "port_a_driver.sv"
`include "port_a_monitor.sv"

endpackage
